library verilog;
use verilog.vl_types.all;
entity DEUARC_group34_vlg_vec_tst is
end DEUARC_group34_vlg_vec_tst;
