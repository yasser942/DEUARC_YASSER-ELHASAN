library verilog;
use verilog.vl_types.all;
entity DEUARC_group34_vlg_check_tst is
    port(
        OutputR         : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end DEUARC_group34_vlg_check_tst;
