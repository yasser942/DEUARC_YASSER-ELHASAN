library verilog;
use verilog.vl_types.all;
entity DEUARC_group34 is
    port(
        OutputR         : out    vl_logic_vector(3 downto 0);
        Clock           : in     vl_logic;
        InputR          : in     vl_logic_vector(3 downto 0)
    );
end DEUARC_group34;
